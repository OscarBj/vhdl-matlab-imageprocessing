-- CCL algorithm